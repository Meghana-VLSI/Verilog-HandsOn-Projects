`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 18.10.2025 18:50:32
// Design Name: 
// Module Name: parallel_adder_4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



// 4-bit Parallel Adder using 4 Full Adders
module parallel_adder_4 (
    input [3:0]a,b,
    input cin,
    output [3:0]sum,
    output cout
);
    wire c1, c2, c3; 
    
    full_adder FA0 (.a(a[0]),.b( b[0]), .cin(cin),.sum( sum[0]),.cout( c1));
    full_adder FA1 (.a(a[1]),.b( b[1]),.cin( c1),.sum(sum[1]),.cout( c2));
    full_adder FA2 (.a(a[2]),.b( b[2]),.cin( c2),.sum(sum[2]),.cout( c3));
    full_adder FA3 (.a(a[3]),.b( b[3]),.cin( c3),.sum( sum[3]),.cout( cout));

endmodule
